/*----------------------------------------------------------------
  Testbench
------------------------------------------------------------------*/
module tb_lab6 ();

logic clk , reset;

Project_1 uut (.clk(clk), .reset(reset));
parameter T = 10; // Clock Period
/*----------------------------------------------------------------
  Clock Generator
------------------------------------------------------------------*/
initial
begin
clk = 0;
forever #(T/2) clk=~clk;
end

initial
begin
reset = 1;
@(posedge clk);
reset = 0;
#110;
end
/*----------------------------------------------------------------
  Reset Sequence
------------------------------------------------------------------*/

endmodule